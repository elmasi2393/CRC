----------------------------------------------------------------------------------
-- Company: Universidad Tecnol�gica Nacional - Facultad Regional San Francisco
-- Engineer: Rinaudo, Facundo. Gatto, Maximiliano. Lenta, Maximiliano.
-- 
-- Create Date:    18:49:34 07/13/2020 
-- Design Name: T�cnicas Digitales I. Trabajo Pr�ctico N�3
-- Module Name:    CRC - COMPORTAMIENTO 
-- Project Name: Dise�o Circuito Generador CRC

-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity CRC is
	GENERIC(M: INTEGER:=8;
				N: INTEGER:=4);
		
		PORT(MENSAJE: IN STD_LOGIC_VECTOR(M-1 DOWNTO 0);	--MENSAJE DE 8 BITS
				POLGEN: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);	--POLINOMIO GENERADOR 4 BITS
				
				BITSCOMP: OUT STD_LOGIC_VECTOR(N-2 DOWNTO 0);	--3 BITS DE COMPROBACI�N
				MENSBITSCOMP: OUT STD_LOGIC_VECTOR(M+N-2 DOWNTO 0));	--8 BITS MENSAJE DE ENTRADA + 3 BITS DE COMPROBACI�N
end CRC;

architecture COMPORTAMIENTO of CRC is

begin
	PROCESS(MENSAJE, POLGEN)
		VARIABLE VAR1: STD_LOGIC_VECTOR(M+N-2 DOWNTO 0); --11 bits - 10 downto 0
		VARIABLE VAR2: STD_LOGIC_VECTOR(N-1 DOWNTO 0); --Variables de 4 bits
		VARIABLE VAR3: STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		VARIABLE VAR4: STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		
	BEGIN
		VAR1(M+N-2 DOWNTO N-1):=MENSAJE(M-1 DOWNTO 0);	--ALMACENA EN LAS POSICIONES (10 DOWNTO 3) DEL VACTOR VAR1
																			--LAS POSICIONES (7 DOWNTO 0) DEL VECTOR MENSAJE
		
		FOR j IN N-2 DOWNTO 0 LOOP		--INICIALIZA LAS POSICIONES (2 DOWNTO 0) DEL VECTOR VAR1 EN CERO
			VAR1(j):='0';
			END LOOP;
			
		VAR2:=POLGEN;	--ALMACENA LOS BITS DEL POLINOMIO GENERADOR EN EL VECTOR VAR2
		
		VAR3:=VAR1(M+N-2 DOWNTO M-1);		--ALMACENA LAS POSICIONES (10 DOWNTO 7) DEL VECTOR VAR1, EN EL VECTOR VAR3
														--ES DECIR, LOS CUATRO BITS MAS SIGNIFICATIVOS EL MENSAJE
		
		FOR i IN M-1 DOWNTO 0 LOOP
			IF(VAR3(N-1)='1') THEN		--ANALIZA SI EL BIT MAS SIGNIFICATIVO DEL VECTOR MENSAJE ES IGUAL A 1
				VAR3:=VAR3 XOR VAR2;			--SI ES AS�, REALIZA LA OPERACI�N XOR ENTRE LAS POSICIONES (3 DOWNTO 0) DE VAR3 
														--Y LAS POSICIONES (3 DOWNTO 0) DEL POLINOMIO GENERADOR. 
				ELSE											--DE LO CONTRARIO VAR3 PERMANECE SIN CAMBIOS
					NULL;
				
			END IF;
		
		VAR4:=VAR3;	--ALMACENA VAR3 EN VAR 4
		
		VAR3(N-1 DOWNTO 1):=VAR4(N-2 DOWNTO 0);	--ALMACENA EN LAS POSICIONES (3 DOWNTO 1) DE VAR3 
																	--LAS POSICIONES (2 DOWNTO 0) DE VAR4 
			IF(i=0) THEN
				VAR3(0):='0';	--SI i=0 ENTONCES ASIGNA CERO A VAR3(0)
				
				ELSE	--DE LO CONTRARIOASIGNA EL VALOR (i-1) A LA POSICI�N VAR3(0)
					VAR3(0):=VAR1(i-1);
				
			END IF;
			
		END LOOP;
		
		BITSCOMP<=VAR3(N-1 DOWNTO 1);	--ASIGNA A BITSCOMP LAS POSICIONES (3 DOWNTO 0) DEL VECTOR VAR3
		
		MENSBITSCOMP(M+N-2 DOWNTO N-1)<=MENSAJE;	--ASIGNA A LAS POSICIONES (10 DOWNTO 3) LOS BITS CORRESPONDIENTES
																	--AL MENSAJE QUE SE DESEA ENVIAR
		MENSBITSCOMP(N-2 DOWNTO 0)<=VAR3(N-1 DOWNTO 1);	--Y A LAS POSICIONES (2 DOWNTO 0) LOS BITS CORRESPONDIENTES
																			--A LAS POSICIONES (3 DOWNTO 1) DE VAR3
	END PROCESS;
														
end COMPORTAMIENTO;

